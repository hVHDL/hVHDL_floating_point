library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package denormalizer_pipeline_pkg is

    constant pipeline_configuration : natural := 1;

end package denormalizer_pipeline_pkg;
