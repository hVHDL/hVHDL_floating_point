LIBRARY ieee  ; 
    USE ieee.NUMERIC_STD.all  ; 
    USE ieee.std_logic_1164.all  ; 
    use ieee.math_real.all;

    use work.float_type_definitions_pkg.all;
    use work.float_arithmetic_operations_pkg.all;
    use work.float_to_real_conversions_pkg.all;

library vunit_lib;
    use vunit_lib.run_pkg.all;

entity float_conversions_tb is
  generic (runner_cfg : string);
end;

architecture vunit_simulation of float_conversions_tb is

    signal simulation_running : boolean;
    signal simulator_clock : std_logic;
    constant clock_per : time := 1 ns;
    constant clock_half_per : time := 0.5 ns;
    constant simtime_in_clocks : integer := 50;

    signal simulation_counter : natural := 0;
    -----------------------------------
    -- simulation specific signals ----
    constant init_test_1 : float_record := to_float(568996.25);
    constant init_test_2 : float_record := to_float(4.0);
    constant init_test_3 : float_record := to_float(-3.2);
    constant init_test_4 : float_record := to_float(8.0);

    signal test_1 : float_record := init_test_1;
    signal test_2 : float_record := init_test_2;
    signal test_3 : float_record := init_test_3;
    signal test_4 : float_record := init_test_4;

    signal test_1_real: real := to_real(init_test_1);
    signal test_2_real: real := to_real(init_test_2);
    signal test_3_real: real := to_real(init_test_3);
    signal test_4_real: real := to_real(init_test_4);

    constant init_test_float : float_record := to_float(22.1346836);
    signal test_float : float_record := init_test_float;
    signal test_real : real := to_real(init_test_float);


------------------------------------------------------------------------

begin

------------------------------------------------------------------------
    simtime : process
    begin
        test_runner_setup(runner, runner_cfg);
        simulation_running <= true;
        wait for simtime_in_clocks*clock_per;
        simulation_running <= false;
        test_runner_cleanup(runner); -- Simulation ends here
        wait;
    end process simtime;	

------------------------------------------------------------------------
    sim_clock_gen : process
    begin
        simulator_clock <= '0';
        wait for clock_half_per;
        while simulation_running loop
            wait for clock_half_per;
                simulator_clock <= not simulator_clock;
            end loop;
        wait;
    end process;
------------------------------------------------------------------------

    stimulus : process(simulator_clock)

    begin
        if rising_edge(simulator_clock) then
            simulation_counter <= simulation_counter + 1;

        end if; -- rising_edge
    end process stimulus;	
------------------------------------------------------------------------
end vunit_simulation;
