library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

    use work.float_type_definitions_pkg.all;

package float_arithmetic_operations_pkg is
    package( package float_typedefs is new work.float_type_definitions_pkg generic map(<>));

end package float_arithmetic_operations_pkg;


package body float_arithmetic_operations_pkg is
end package body float_arithmetic_operations_pkg;
