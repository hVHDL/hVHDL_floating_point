library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;


-- 24 bits
package float_word_length_pkg is

    constant mantissa_bits : integer := 24;
    constant exponent_bits : integer := 8;

end package float_word_length_pkg;

