library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

    use work.float_type_definitions_pkg.all;
    use work.float_adder_pkg.all;
    use work.float_multiplier_pkg.all;
    use work.normalizer_pkg.all;

package float_alu_pkg is
------------------------------------------------------------------------
    type float_alu_record is record

        float_adder                 : float_adder_record      ;
        float_adder_normalizer      : float_normalizer_record ;

        float_multiplier            : float_multiplier_record ;
        float_multiplier_normalizer : float_normalizer_record ;

        float_alu_is_busy : boolean;
    end record;

    constant init_float_alu : float_alu_record := (
            init_float_adder      ,
            init_float_normalizer ,

            init_float_multiplier ,
            init_float_normalizer ,

            false);

------------------------------------------------------------------------
    procedure create_float_alu (
        signal float_alu_object : inout float_alu_record);
------------------------------------------------------------------------
end package float_alu_pkg;

package body float_alu_pkg is
------------------------------------------------------------------------
    procedure create_float_alu 
    (
        signal float_alu_object : inout float_alu_record
    ) 
    is

        alias float_adder                 is float_alu_object.float_adder                ;
        alias float_multiplier            is float_alu_object.float_multiplier           ;
        alias float_adder_normalizer      is float_alu_object.float_adder_normalizer     ;
        alias float_multiplier_normalizer is float_alu_object.float_multiplier_normalizer;
    begin

        create_adder(float_adder);
        create_normalizer(float_adder_normalizer);

        create_float_multiplier(float_multiplier);
        create_normalizer(float_multiplier_normalizer);

    end procedure;
------------------------------------------------------------------------
------------------------------------------------------------------------
    procedure multiply
    (
        signal alu_object : inout float_alu_record;
        left, right : float_record
    ) is
    begin

        request_float_multiplier(
            alu_object.float_multiplier,
            left, right);
    end multiply;
------------------------------------------------------------------------
    function multiplier_is_ready
    (
        alu_object : float_alu_record
    )
    return boolean
    is
    begin
        return float_multiplier_is_ready(alu_object.float_multiplier);
    end multiplier_is_ready;
------------------------------------------------------------------------
    function get_multiplier_result
    (
        alu_object : float_alu_record
    )
    return float_record
    is
    begin
        return get_multiplier_result(alu_object.float_multiplier);
    end get_multiplier_result;
------------------------------------------------------------------------
------------------------------------------------------------------------
    procedure add
    (
        signal alu_object : inout float_alu_record;
        left, right : float_record
    ) is
    begin
        request_add(alu_object.float_adder, left, right);
    end add;
------------------------------------------------------------------------
end package body float_alu_pkg;
